--------------------------------------------------------------------------------
-- VGA MOTOR
-- Anders Nilsson
-- 16-feb-2016
-- Version 1.1


-- library declaration
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;            -- basic IEEE library
use IEEE.NUMERIC_STD.ALL;               -- IEEE library for the unsigned type


-- entity
entity VGA_MOTOR is
    port ( clk	  : in std_logic;
    	 addr     : out unsigned(12 downto 0);
    	 rst      : in std_logic;
    	 vgaRed   : out std_logic_vector(2 downto 0);
    	 vgaGreen : out std_logic_vector(2 downto 0);
    	 vgaBlue  : out std_logic_vector(2 downto 1);
    	 Hsync    : out std_logic;
    	 Vsync    : out std_logic;
         picmem_in      : in std_logic_vector(7 downto 0);      -- data
         bitmem_in      : in std_logic;      -- data
         Xpixel   : buffer unsigned(9 downto 0);         -- Horizontal pixel counter
         Ypixel   : buffer unsigned(9 downto 0)
         );
end VGA_MOTOR;


-- architecture
architecture Behavioral of VGA_MOTOR is


    signal ClkDiv : unsigned(1 downto 0);		-- Clock divisor, to generate 25 MHz signal
    signal Clk25  : std_logic;			-- One pulse width 25 MHz signal

    signal tilePixel : std_logic_vector(7 downto 0);	-- Tile pixel data
    signal tileAddr  : unsigned(14 downto 0);	-- Tile address

    signal blank : std_logic;                    -- blanking signal
    signal tilerow : std_logic;

    -- Tile memory type
    type ram_t is array (0 to 6143) of std_logic;

signal tileMem : ram_t :=(
        -- 0
        '0','0','0','0','0','0','0','0',
        '0','0','0','0','0','0','0','0',
        '0','0','0','0','0','0','0','0',
        '0','0','0','1','1','0','0','0',
        '0','0','1','0','0','1','0','0',
        '0','1','0','0','0','0','1','0',
        '0','1','0','0','0','0','1','0',
        '0','1','0','1','1','0','1','0',
        '0','1','0','1','1','0','1','0',
        '0','1','0','0','0','0','1','0',
        '0','1','0','0','0','0','1','0',
        '0','0','1','0','0','1','0','0',
        '0','0','0','1','1','0','0','0',
        '0','0','0','0','0','0','0','0',
        '0','0','0','0','0','0','0','0',
        '0','0','0','0','0','0','0','0',
        -- 1
        '0','0','0','0','0','0','0','0',
        '0','0','0','0','0','0','0','0',
        '0','0','0','0','0','0','0','0',
        '0','0','0','0','0','1','0','0',
        '0','0','0','0','1','1','0','0',
        '0','0','0','1','0','1','0','0',
        '0','0','0','0','0','1','0','0',
        '0','0','0','0','0','1','0','0',
        '0','0','0','0','0','1','0','0',
        '0','0','0','0','0','1','0','0',
        '0','0','0','0','0','1','0','0',
        '0','0','0','0','0','1','0','0',
        '0','0','0','1','1','1','1','1',
        '0','0','0','0','0','0','0','0',
        '0','0','0','0','0','0','0','0',
        '0','0','0','0','0','0','0','0',
        -- 2
        '0','0','0','0','0','0','0','0',
        '0','0','0','0','0','0','0','0',
        '0','0','0','0','0','0','0','0',
        '0','0','1','1','1','1','0','0',
        '0','1','0','0','0','0','1','0',
        '0','0','0','0','0','0','1','0',
        '0','0','0','0','0','0','1','0',
        '0','0','0','0','0','1','0','0',
        '0','0','0','0','1','0','0','0',
        '0','0','0','1','0','0','0','0',
        '0','0','1','0','0','0','0','0',
        '0','1','0','0','0','0','0','0',
        '0','1','1','1','1','1','1','0',
        '0','0','0','0','0','0','0','0',
        '0','0','0','0','0','0','0','0',
        '0','0','0','0','0','0','0','0',
        -- 3
        '0','0','0','0','0','0','0','0',
        '0','0','0','0','0','0','0','0',
        '0','0','0','0','0','0','0','0',
        '0','1','1','1','1','1','0','0',
        '0','0','0','0','0','0','1','0',
        '0','0','0','0','0','0','1','0',
        '0','0','0','0','0','0','1','0',
        '0','0','0','1','1','1','0','0',
        '0','0','0','0','0','0','1','0',
        '0','0','0','0','0','0','1','0',
        '0','0','0','0','0','0','1','0',
        '0','0','0','0','0','0','1','0',
        '0','1','1','1','1','1','0','0',
        '0','0','0','0','0','0','0','0',
        '0','0','0','0','0','0','0','0',
        '0','0','0','0','0','0','0','0',
        -- 4
        '0','0','0','0','0','0','0','0',
        '0','0','0','0','0','0','0','0',
        '0','0','0','0','0','0','0','0',
        '0','0','0','0','0','1','0','0',
        '0','0','0','0','1','1','0','0',
        '0','0','0','1','0','1','0','0',
        '0','0','1','0','0','1','0','0',
        '0','0','1','0','0','1','0','0',
        '0','1','0','0','0','1','0','0',
        '0','1','1','1','1','1','1','0',
        '0','0','0','0','0','1','0','0',
        '0','0','0','0','0','1','0','0',
        '0','0','0','0','0','1','0','0',
        '0','0','0','0','0','0','0','0',
        '0','0','0','0','0','0','0','0',
        '0','0','0','0','0','0','0','0',
        -- 5
        '0','0','0','0','0','0','0','0',
        '0','0','0','0','0','0','0','0',
        '0','0','0','0','0','0','0','0',
        '0','0','0','1','1','1','1','1',
        '0','0','0','1','0','0','0','0',
        '0','0','0','1','0','0','0','0',
        '0','0','0','1','0','0','0','0',
        '0','0','0','1','1','1','0','0',
        '0','0','0','0','0','0','1','0',
        '0','0','0','0','0','0','0','1',
        '0','0','0','0','0','0','0','1',
        '0','0','0','0','0','0','1','0',
        '0','0','1','1','1','1','0','0',
        '0','0','0','0','0','0','0','0',
        '0','0','0','0','0','0','0','0',
        '0','0','0','0','0','0','0','0',
        -- 6
        '0','0','0','0','0','0','0','0',
        '0','0','0','0','0','0','0','0',
        '0','0','0','0','0','0','0','0',
        '0','0','0','0','1','1','0','0',
        '0','0','0','1','0','0','0','0',
        '0','0','1','0','0','0','0','0',
        '0','1','0','0','0','0','0','0',
        '0','1','1','1','1','1','0','0',
        '0','1','0','0','0','0','1','0',
        '0','1','0','0','0','0','1','0',
        '0','1','0','0','0','0','1','0',
        '0','0','1','0','0','1','0','0',
        '0','0','0','1','1','0','0','0',
        '0','0','0','0','0','0','0','0',
        '0','0','0','0','0','0','0','0',
        '0','0','0','0','0','0','0','0',
        -- 7
        '0','0','0','0','0','0','0','0',
        '0','0','0','0','0','0','0','0',
        '0','0','0','0','0','0','0','0',
        '0','0','1','1','1','1','1','1',
        '0','0','0','0','0','0','0','1',
        '0','0','0','0','0','0','1','0',
        '0','0','0','0','0','1','0','0',
        '0','0','0','0','0','1','0','0',
        '0','0','0','0','1','0','0','0',
        '0','0','0','0','1','0','0','0',
        '0','0','0','1','0','0','0','0',
        '0','0','0','1','0','0','0','0',
        '0','0','0','1','0','0','0','0',
        '0','0','0','0','0','0','0','0',
        '0','0','0','0','0','0','0','0',
        '0','0','0','0','0','0','0','0',
        -- 8
        '0','0','0','0','0','0','0','0',
        '0','0','0','0','0','0','0','0',
        '0','0','0','0','0','0','0','0',
        '0','0','1','1','1','1','0','0',
        '0','1','0','0','0','0','1','0',
        '0','1','0','0','0','0','1','0',
        '0','1','0','0','0','0','1','0',
        '0','0','1','1','1','1','0','0',
        '0','0','1','0','1','1','0','0',
        '0','1','0','0','0','0','1','0',
        '0','1','0','0','0','0','1','0',
        '0','1','0','0','0','0','1','0',
        '0','0','1','1','1','1','0','0',
        '0','0','0','0','0','0','0','0',
        '0','0','0','0','0','0','0','0',
        '0','0','0','0','0','0','0','0',
        -- 9
        '0','0','0','0','0','0','0','0',
        '0','0','0','0','0','0','0','0',
        '0','0','0','0','0','0','0','0',
        '0','0','1','1','1','0','0','0',
        '0','1','0','0','0','1','0','0',
        '0','1','0','0','0','0','1','0',
        '0','1','0','0','0','0','1','0',
        '0','1','0','0','0','0','1','0',
        '0','0','1','1','1','1','1','0',
        '0','0','0','0','0','0','1','0',
        '0','0','0','0','0','1','0','0',
        '0','0','0','0','1','0','0','0',
        '0','0','1','1','0','0','0','0',
        '0','0','0','0','0','0','0','0',
        '0','0','0','0','0','0','0','0',
        '0','0','0','0','0','0','0','0',
        -- A
        '0','0','0','0','0','0','0','0',
        '0','0','0','0','0','0','0','0',
        '0','0','0','0','0','0','0','0',
        '0','0','0','1','0','0','0','0',
        '0','0','1','0','1','0','0','0',
        '0','0','1','0','1','0','0','0',
        '0','0','1','0','1','0','0','0',
        '0','1','0','0','0','1','0','0',
        '0','1','0','0','0','1','0','0',
        '0','1','1','1','1','1','0','0',
        '0','1','0','0','0','1','0','0',
        '1','0','0','0','0','0','1','0',
        '1','0','0','0','0','0','1','0',
        '0','0','0','0','0','0','0','0',
        '0','0','0','0','0','0','0','0',
        '0','0','0','0','0','0','0','0',
        -- B
        '0','0','0','0','0','0','0','0',
        '0','0','0','0','0','0','0','0',
        '0','0','0','0','0','0','0','0',
        '0','1','1','1','1','1','0','0',
        '0','1','0','0','0','0','1','0',
        '0','1','0','0','0','0','1','0',
        '0','1','0','0','0','0','1','0',
        '0','1','1','1','1','1','0','0',
        '0','1','0','0','0','0','1','0',
        '0','1','0','0','0','0','1','0',
        '0','1','0','0','0','0','1','0',
        '0','1','0','0','0','0','1','0',
        '0','1','1','1','1','1','0','0',
        '0','0','0','0','0','0','0','0',
        '0','0','0','0','0','0','0','0',
        '0','0','0','0','0','0','0','0',
        -- C
        '0','0','0','0','0','0','0','0',
        '0','0','0','0','0','0','0','0',
        '0','0','0','0','0','0','0','0',
        '0','0','0','1','1','1','0','0',
        '0','0','1','0','0','0','1','0',
        '0','1','0','0','0','0','0','0',
        '0','1','0','0','0','0','0','0',
        '0','1','0','0','0','0','0','0',
        '0','1','0','0','0','0','0','0',
        '0','1','0','0','0','0','0','0',
        '0','1','0','0','0','0','0','0',
        '0','0','1','0','0','0','1','0',
        '0','0','0','1','1','1','0','0',
        '0','0','0','0','0','0','0','0',
        '0','0','0','0','0','0','0','0',
        '0','0','0','0','0','0','0','0',
        -- D
        '0','0','0','0','0','0','0','0',
        '0','0','0','0','0','0','0','0',
        '0','0','0','0','0','0','0','0',
        '0','1','1','1','1','0','0','0',
        '0','1','0','0','0','1','0','0',
        '0','1','0','0','0','0','1','0',
        '0','1','0','0','0','0','1','0',
        '0','1','0','0','0','0','1','0',
        '0','1','0','0','0','0','1','0',
        '0','1','0','0','0','0','1','0',
        '0','1','0','0','0','0','1','0',
        '0','1','0','0','0','1','0','0',
        '0','1','1','1','1','0','0','0',
        '0','0','0','0','0','0','0','0',
        '0','0','0','0','0','0','0','0',
        '0','0','0','0','0','0','0','0',
        -- E
        '0','0','0','0','0','0','0','0',
        '0','0','0','0','0','0','0','0',
        '0','0','0','0','0','0','0','0',
        '0','0','1','1','1','1','1','1',
        '0','0','1','0','0','0','0','0',
        '0','0','1','0','0','0','0','0',
        '0','0','1','0','0','0','0','0',
        '0','0','1','1','1','1','1','0',
        '0','0','1','0','0','0','0','0',
        '0','0','1','0','0','0','0','0',
        '0','0','1','0','0','0','0','0',
        '0','0','1','0','0','0','0','0',
        '0','0','1','1','1','1','1','1',
        '0','0','0','0','0','0','0','0',
        '0','0','0','0','0','0','0','0',
        '0','0','0','0','0','0','0','0',
        -- F
        '0','0','0','0','0','0','0','0',
        '0','0','0','0','0','0','0','0',
        '0','0','0','0','0','0','0','0',
        '0','0','1','1','1','1','1','1',
        '0','0','1','0','0','0','0','0',
        '0','0','1','0','0','0','0','0',
        '0','0','1','0','0','0','0','0',
        '0','0','1','1','1','1','1','0',
        '0','0','1','0','0','0','0','0',
        '0','0','1','0','0','0','0','0',
        '0','0','1','0','0','0','0','0',
        '0','0','1','0','0','0','0','0',
        '0','0','1','0','0','0','0','0',
        '0','0','0','0','0','0','0','0',
        '0','0','0','0','0','0','0','0',
        '0','0','0','0','0','0','0','0',
        -- G
        '0','0','0','0','0','0','0','0',
        '0','0','0','0','0','0','0','0',
        '0','0','0','0','0','0','0','0',
        '0','0','0','1','1','1','0','0',
        '0','0','1','0','0','0','1','0',
        '0','1','0','0','0','0','0','0',
        '0','1','0','0','0','0','0','0',
        '0','1','0','0','0','0','0','0',
        '0','1','0','0','0','0','1','0',
        '0','1','0','0','0','0','1','0',
        '0','1','0','0','0','0','1','0',
        '0','0','1','0','0','0','1','0',
        '0','0','0','1','1','1','1','0',
        '0','0','0','0','0','0','0','0',
        '0','0','0','0','0','0','0','0',
        '0','0','0','0','0','0','0','0',
        -- H
        '0','0','0','0','0','0','0','0',
        '0','0','0','0','0','0','0','0',
        '0','0','0','0','0','0','0','0',
        '0','1','0','0','0','0','1','0',
        '0','1','0','0','0','0','1','0',
        '0','1','0','0','0','0','1','0',
        '0','1','0','0','0','0','1','0',
        '0','1','1','1','1','1','1','0',
        '0','1','0','0','0','0','1','0',
        '0','1','0','0','0','0','1','0',
        '0','1','0','0','0','0','1','0',
        '0','1','0','0','0','0','1','0',
        '0','1','0','0','0','0','1','0',
        '0','0','0','0','0','0','0','0',
        '0','0','0','0','0','0','0','0',
        '0','0','0','0','0','0','0','0',
        -- I
        '0','0','0','0','0','0','0','0',
        '0','0','0','0','0','0','0','0',
        '0','0','0','0','0','0','0','0',
        '0','0','1','1','1','1','1','0',
        '0','0','0','0','1','0','0','0',
        '0','0','0','0','1','0','0','0',
        '0','0','0','0','1','0','0','0',
        '0','0','0','0','1','0','0','0',
        '0','0','0','0','1','0','0','0',
        '0','0','0','0','1','0','0','0',
        '0','0','0','0','1','0','0','0',
        '0','0','0','0','1','0','0','0',
        '0','0','1','1','1','1','1','0',
        '0','0','0','0','0','0','0','0',
        '0','0','0','0','0','0','0','0',
        '0','0','0','0','0','0','0','0',
        -- J
        '0','0','0','0','0','0','0','0',
        '0','0','0','0','0','0','0','0',
        '0','0','0','0','0','0','0','0',
        '0','0','1','1','1','1','1','0',
        '0','0','0','0','0','0','1','0',
        '0','0','0','0','0','0','1','0',
        '0','0','0','0','0','0','1','0',
        '0','0','0','0','0','0','1','0',
        '0','0','0','0','0','0','1','0',
        '0','0','0','0','0','0','1','0',
        '0','0','0','0','0','0','1','0',
        '0','1','0','0','0','0','1','0',
        '0','0','1','1','1','1','0','0',
        '0','0','0','0','0','0','0','0',
        '0','0','0','0','0','0','0','0',
        '0','0','0','0','0','0','0','0',
        -- K
        '0','0','0','0','0','0','0','0',
        '0','0','0','0','0','0','0','0',
        '0','0','0','0','0','0','0','0',
        '0','0','1','0','0','0','0','1',
        '0','0','1','0','0','0','1','0',
        '0','0','1','0','0','1','0','0',
        '0','0','1','0','1','0','0','0',
        '0','0','1','1','0','0','0','0',
        '0','0','1','0','1','0','0','0',
        '0','0','1','0','0','1','0','0',
        '0','0','1','0','0','1','0','0',
        '0','0','1','0','0','0','1','0',
        '0','0','1','0','0','0','0','1',
        '0','0','0','0','0','0','0','0',
        '0','0','0','0','0','0','0','0',
        '0','0','0','0','0','0','0','0',
        -- L
        '0','0','0','0','0','0','0','0',
        '0','0','0','0','0','0','0','0',
        '0','0','0','0','0','0','0','0',
        '0','0','1','0','0','0','0','0',
        '0','0','1','0','0','0','0','0',
        '0','0','1','0','0','0','0','0',
        '0','0','1','0','0','0','0','0',
        '0','0','1','0','0','0','0','0',
        '0','0','1','0','0','0','0','0',
        '0','0','1','0','0','0','0','0',
        '0','0','1','0','0','0','0','0',
        '0','0','1','0','0','0','0','0',
        '0','0','1','1','1','1','1','1',
        '0','0','0','0','0','0','0','0',
        '0','0','0','0','0','0','0','0',
        '0','0','0','0','0','0','0','0',
        -- M
        '0','0','0','0','0','0','0','0',
        '0','0','0','0','0','0','0','0',
        '0','0','0','0','0','0','0','0',
        '0','0','1','0','0','1','0','0',
        '0','0','1','0','0','1','0','0',
        '0','0','1','0','0','1','0','0',
        '0','1','0','1','1','0','1','0',
        '0','1','0','1','1','0','1','0',
        '0','1','0','1','1','0','1','0',
        '0','1','0','0','0','0','1','0',
        '0','1','0','0','0','0','1','0',
        '0','1','0','0','0','0','1','0',
        '0','1','0','0','0','0','1','0',
        '0','0','0','0','0','0','0','0',
        '0','0','0','0','0','0','0','0',
        '0','0','0','0','0','0','0','0',
        -- N
        '0','0','0','0','0','0','0','0',
        '0','0','0','0','0','0','0','0',
        '0','0','0','0','0','0','0','0',
        '0','1','0','0','0','0','1','0',
        '0','1','1','0','0','0','1','0',
        '0','1','1','0','0','0','1','0',
        '0','1','0','1','0','0','1','0',
        '0','1','0','1','1','0','1','0',
        '0','1','0','0','1','0','1','0',
        '0','1','0','0','1','0','1','0',
        '0','1','0','0','0','1','1','0',
        '0','1','0','0','0','1','1','0',
        '0','1','0','0','0','0','1','0',
        '0','0','0','0','0','0','0','0',
        '0','0','0','0','0','0','0','0',
        '0','0','0','0','0','0','0','0',
        -- O
        '0','0','0','0','0','0','0','0',
        '0','0','0','0','0','0','0','0',
        '0','0','0','0','0','0','0','0',
        '0','0','0','1','1','0','0','0',
        '0','0','1','0','0','1','0','0',
        '0','1','0','0','0','0','1','0',
        '0','1','0','0','0','0','1','0',
        '0','1','0','0','0','0','1','0',
        '0','1','0','0','0','0','1','0',
        '0','1','0','0','0','0','1','0',
        '0','1','0','0','0','0','1','0',
        '0','0','1','0','0','1','0','0',
        '0','0','0','1','1','0','0','0',
        '0','0','0','0','0','0','0','0',
        '0','0','0','0','0','0','0','0',
        '0','0','0','0','0','0','0','0',
        -- P
        '0','0','0','0','0','0','0','0',
        '0','0','0','0','0','0','0','0',
        '0','0','0','0','0','0','0','0',
        '0','0','1','1','1','1','1','0',
        '0','0','1','0','0','0','0','1',
        '0','0','1','0','0','0','0','1',
        '0','0','1','0','0','0','0','1',
        '0','0','1','0','0','0','0','1',
        '0','0','1','1','1','1','1','0',
        '0','0','1','0','0','0','0','0',
        '0','0','1','0','0','0','0','0',
        '0','0','1','0','0','0','0','0',
        '0','0','1','0','0','0','0','0',
        '0','0','0','0','0','0','0','0',
        '0','0','0','0','0','0','0','0',
        '0','0','0','0','0','0','0','0',
        -- Q
        '0','0','0','0','0','0','0','0',
        '0','0','0','0','0','0','0','0',
        '0','0','0','0','0','0','0','0',
        '0','0','0','1','1','0','0','0',
        '0','0','1','0','0','1','0','0',
        '0','1','0','0','0','0','1','0',
        '0','1','0','0','0','0','1','0',
        '0','1','0','0','0','0','1','0',
        '0','1','0','0','0','0','1','0',
        '0','1','0','0','0','0','1','0',
        '0','1','0','0','0','0','1','0',
        '0','0','1','0','0','1','0','0',
        '0','0','0','1','1','0','0','0',
        '0','0','0','1','1','0','0','0',
        '0','0','0','0','0','1','1','0',
        '0','0','0','0','0','0','0','0',
        -- R
        '0','0','0','0','0','0','0','0',
        '0','0','0','0','0','0','0','0',
        '0','0','0','0','0','0','0','0',
        '0','1','1','1','1','1','0','0',
        '0','1','0','0','0','0','1','0',
        '0','1','0','0','0','0','1','0',
        '0','1','0','0','0','0','1','0',
        '0','1','0','0','0','0','1','0',
        '0','1','1','1','1','1','0','0',
        '0','1','0','0','1','0','0','0',
        '0','1','0','0','0','1','0','0',
        '0','1','0','0','0','0','1','0',
        '0','1','0','0','0','0','0','1',
        '0','0','0','0','0','0','0','0',
        '0','0','0','0','0','0','0','0',
        '0','0','0','0','0','0','0','0',
        -- S
        '0','0','0','0','0','0','0','0',
        '0','0','0','0','0','0','0','0',
        '0','0','0','0','0','0','0','0',
        '0','0','1','1','1','1','0','0',
        '0','1','0','0','0','0','1','0',
        '0','1','0','0','0','0','0','0',
        '0','1','0','0','0','0','0','0',
        '0','0','1','1','0','0','0','0',
        '0','0','0','0','1','1','0','0',
        '0','0','0','0','0','0','1','0',
        '0','0','0','0','0','0','1','0',
        '0','1','0','0','0','0','1','0',
        '0','1','1','1','1','1','0','0',
        '0','0','0','0','0','0','0','0',
        '0','0','0','0','0','0','0','0',
        '0','0','0','0','0','0','0','0',
        -- T
        '0','0','0','0','0','0','0','0',
        '0','0','0','0','0','0','0','0',
        '0','0','0','0','0','0','0','0',
        '1','1','1','1','1','1','1','0',
        '0','0','0','1','0','0','0','0',
        '0','0','0','1','0','0','0','0',
        '0','0','0','1','0','0','0','0',
        '0','0','0','1','0','0','0','0',
        '0','0','0','1','0','0','0','0',
        '0','0','0','1','0','0','0','0',
        '0','0','0','1','0','0','0','0',
        '0','0','0','1','0','0','0','0',
        '0','0','0','1','0','0','0','0',
        '0','0','0','0','0','0','0','0',
        '0','0','0','0','0','0','0','0',
        '0','0','0','0','0','0','0','0',
        -- U
        '0','0','0','0','0','0','0','0',
        '0','0','0','0','0','0','0','0',
        '0','0','0','0','0','0','0','0',
        '0','1','0','0','0','0','1','0',
        '0','1','0','0','0','0','1','0',
        '0','1','0','0','0','0','1','0',
        '0','1','0','0','0','0','1','0',
        '0','1','0','0','0','0','1','0',
        '0','1','0','0','0','0','1','0',
        '0','1','0','0','0','0','1','0',
        '0','1','0','0','0','0','1','0',
        '0','1','0','0','0','0','1','0',
        '0','0','1','1','1','1','0','0',
        '0','0','0','0','0','0','0','0',
        '0','0','0','0','0','0','0','0',
        '0','0','0','0','0','0','0','0',
        -- V
        '0','0','0','0','0','0','0','0',
        '0','0','0','0','0','0','0','0',
        '0','0','0','0','0','0','0','0',
        '1','0','0','0','0','0','1','0',
        '1','0','0','0','0','0','1','0',
        '0','1','0','0','0','1','0','0',
        '0','1','0','0','0','1','0','0',
        '0','1','0','0','0','1','0','0',
        '0','1','1','0','0','1','0','0',
        '0','0','1','0','1','0','0','0',
        '0','0','1','0','1','0','0','0',
        '0','0','1','1','1','0','0','0',
        '0','0','0','1','0','0','0','0',
        '0','0','0','0','0','0','0','0',
        '0','0','0','0','0','0','0','0',
        '0','0','0','0','0','0','0','0',
        -- W
        '0','0','0','0','0','0','0','0',
        '0','0','0','0','0','0','0','0',
        '0','0','0','0','0','0','0','0',
        '0','1','0','0','0','0','1','0',
        '0','1','0','0','0','0','1','0',
        '0','1','0','0','0','0','1','0',
        '0','1','0','0','0','0','1','0',
        '0','1','0','1','1','0','1','0',
        '0','1','0','1','1','0','1','0',
        '0','1','0','1','1','0','1','0',
        '0','1','1','0','0','1','1','0',
        '0','1','1','0','0','1','1','0',
        '0','1','0','0','0','0','1','0',
        '0','0','0','0','0','0','0','0',
        '0','0','0','0','0','0','0','0',
        '0','0','0','0','0','0','0','0',
        -- X
        '0','0','0','0','0','0','0','0',
        '0','0','0','0','0','0','0','0',
        '0','0','0','0','0','0','0','0',
        '0','1','0','0','0','0','0','1',
        '0','0','1','0','0','0','1','0',
        '0','0','1','0','0','0','1','0',
        '0','0','0','1','0','1','0','0',
        '0','0','0','0','1','0','0','0',
        '0','0','0','0','1','0','0','0',
        '0','0','0','1','0','1','0','0',
        '0','0','1','0','0','0','1','0',
        '0','0','1','0','0','0','1','0',
        '0','1','0','0','0','0','0','1',
        '0','0','0','0','0','0','0','0',
        '0','0','0','0','0','0','0','0',
        '0','0','0','0','0','0','0','0',
        -- Y
        '0','0','0','0','0','0','0','0',
        '0','0','0','0','0','0','0','0',
        '0','0','0','0','0','0','0','0',
        '1','0','0','0','0','0','1','0',
        '0','1','0','0','0','1','0','0',
        '0','1','0','0','0','1','0','0',
        '0','0','1','0','1','0','0','0',
        '0','0','1','0','1','0','0','0',
        '0','0','0','1','0','0','0','0',
        '0','0','0','1','0','0','0','0',
        '0','0','0','1','0','0','0','0',
        '0','0','0','1','0','0','0','0',
        '0','0','0','1','0','0','0','0',
        '0','0','0','0','0','0','0','0',
        '0','0','0','0','0','0','0','0',
        '0','0','0','0','0','0','0','0',
        -- Z
        '0','0','0','0','0','0','0','0',
        '0','0','0','0','0','0','0','0',
        '0','0','0','0','0','0','0','0',
        '0','1','1','1','1','1','1','0',
        '0','0','0','0','0','0','1','0',
        '0','0','0','0','0','1','0','0',
        '0','0','0','0','1','0','0','0',
        '0','0','0','0','1','0','0','0',
        '0','0','0','1','0','0','0','0',
        '0','0','1','1','0','0','0','0',
        '0','0','1','0','0','0','0','0',
        '0','1','0','0','0','0','0','0',
        '0','1','1','1','1','1','1','0',
        '0','0','0','0','0','0','0','0',
        '0','0','0','0','0','0','0','0',
        '0','0','0','0','0','0','0','0',
        -- Å
        '0','0','0','1','1','0','0','0',
        '0','0','1','0','0','1','0','0',
        '0','0','1','0','0','1','0','0',
        '0','0','0','1','1','0','0','0',
        '0','0','0','1','1','0','0','0',
        '0','0','1','0','0','1','0','0',
        '0','0','1','0','0','1','0','0',
        '0','0','1','0','0','1','0','0',
        '0','1','0','0','0','0','1','0',
        '0','1','1','1','1','1','1','0',
        '0','1','0','0','0','0','1','0',
        '1','0','0','0','0','0','1','1',
        '1','0','0','0','0','0','0','1',
        '0','0','0','0','0','0','0','0',
        '0','0','0','0','0','0','0','0',
        '0','0','0','0','0','0','0','0',
        -- Ä
        '0','0','1','0','1','0','0','0',
        '0','0','1','0','1','0','0','0',
        '0','0','0','0','0','0','0','0',
        '0','0','0','1','0','0','0','0',
        '0','0','1','0','1','0','0','0',
        '0','0','1','0','1','0','0','0',
        '0','0','1','0','1','0','0','0',
        '0','1','0','0','0','1','0','0',
        '0','1','0','0','0','1','0','0',
        '0','1','1','1','1','1','0','0',
        '0','1','0','0','0','1','0','0',
        '1','0','0','0','0','0','1','0',
        '1','0','0','0','0','0','1','0',
        '0','0','0','0','0','0','0','0',
        '0','0','0','0','0','0','0','0',
        '0','0','0','0','0','0','0','0',
        -- Ö
        '0','0','0','1','0','1','0','0',
        '0','0','0','1','0','1','0','0',
        '0','0','0','0','0','0','0','0',
        '0','0','0','1','1','0','0','0',
        '0','0','1','0','0','1','0','0',
        '0','1','0','0','0','0','1','0',
        '0','1','0','0','0','0','1','0',
        '0','1','0','0','0','0','1','0',
        '0','1','0','0','0','0','1','0',
        '0','1','0','0','0','0','1','0',
        '0','1','0','0','0','0','1','0',
        '0','0','1','0','0','1','0','0',
        '0','0','0','1','1','0','0','0',
        '0','0','0','0','0','0','0','0',
        '0','0','0','0','0','0','0','0',
        '0','0','0','0','0','0','0','0',
        -- π
        '0','0','0','0','0','0','0','0',
        '0','0','0','0','0','0','0','0',
        '0','0','0','0','0','0','0','0',
        '0','0','0','0','0','0','0','0',
        '0','0','0','0','0','0','0','0',
        '0','0','0','0','0','0','0','0',
        '0','0','1','1','1','1','1','1',
        '0','0','1','0','0','0','0','1',
        '0','0','1','0','0','0','0','1',
        '0','0','1','0','0','0','0','1',
        '0','0','1','0','0','0','0','1',
        '0','0','1','0','0','0','0','1',
        '0','0','1','0','0','0','0','1',
        '0','0','0','0','0','0','0','0',
        '0','0','0','0','0','0','0','0',
        '0','0','0','0','0','0','0','0',
        -- Ω
        '0','0','0','0','0','0','0','0',
        '0','0','0','0','0','0','0','0',
        '0','0','0','0','0','0','0','0',
        '0','0','0','1','1','0','0','0',
        '0','0','1','0','0','1','0','0',
        '0','1','0','0','0','0','1','0',
        '0','1','0','0','0','0','1','0',
        '0','1','0','0','0','0','1','0',
        '0','1','0','0','0','0','1','0',
        '0','1','0','0','0','0','1','0',
        '0','1','0','0','0','0','1','0',
        '0','0','1','0','0','1','0','0',
        '0','1','1','0','0','1','1','0',
        '0','0','0','0','0','0','0','0',
        '0','0','0','0','0','0','0','0',
        '0','0','0','0','0','0','0','0',
        -- .
        '0','0','0','0','0','0','0','0',
        '0','0','0','0','0','0','0','0',
        '0','0','0','0','0','0','0','0',
        '0','0','0','0','0','0','0','0',
        '0','0','0','0','0','0','0','0',
        '0','0','0','0','0','0','0','0',
        '0','0','0','0','0','0','0','0',
        '0','0','0','0','0','0','0','0',
        '0','0','0','0','0','0','0','0',
        '0','0','0','0','0','0','0','0',
        '0','0','0','0','0','0','0','0',
        '0','0','0','0','0','0','0','0',
        '0','0','0','0','1','0','0','0',
        '0','0','0','0','0','0','0','0',
        '0','0','0','0','0','0','0','0',
        '0','0','0','0','0','0','0','0',
        -- =
        '0','0','0','0','0','0','0','0',
        '0','0','0','0','0','0','0','0',
        '0','0','0','0','0','0','0','0',
        '0','0','0','0','0','0','0','0',
        '0','0','0','0','0','0','0','0',
        '0','0','0','0','0','0','0','0',
        '0','0','0','0','0','0','0','0',
        '0','1','1','1','1','1','1','0',
        '0','0','0','0','0','0','0','0',
        '0','0','0','0','0','0','0','0',
        '0','1','1','1','1','1','1','0',
        '0','0','0','0','0','0','0','0',
        '0','0','0','0','0','0','0','0',
        '0','0','0','0','0','0','0','0',
        '0','0','0','0','0','0','0','0',
        '0','0','0','0','0','0','0','0',
        -- +
        '0','0','0','0','0','0','0','0',
        '0','0','0','0','0','0','0','0',
        '0','0','0','0','0','0','0','0',
        '0','0','0','0','0','0','0','0',
        '0','0','0','0','0','0','0','0',
        '0','0','0','1','0','0','0','0',
        '0','0','0','1','0','0','0','0',
        '0','0','0','1','0','0','0','0',
        '1','1','1','1','1','1','1','0',
        '0','0','0','1','0','0','0','0',
        '0','0','0','1','0','0','0','0',
        '0','0','0','1','0','0','0','0',
        '0','0','0','0','0','0','0','0',
        '0','0','0','0','0','0','0','0',
        '0','0','0','0','0','0','0','0',
        '0','0','0','0','0','0','0','0',
        -- -
        '0','0','0','0','0','0','0','0',
        '0','0','0','0','0','0','0','0',
        '0','0','0','0','0','0','0','0',
        '0','0','0','0','0','0','0','0',
        '0','0','0','0','0','0','0','0',
        '0','0','0','0','0','0','0','0',
        '0','0','0','0','0','0','0','0',
        '0','0','0','0','0','0','0','0',
        '0','0','0','0','0','0','0','0',
        '0','0','0','1','1','1','1','0',
        '0','0','0','0','0','0','0','0',
        '0','0','0','0','0','0','0','0',
        '0','0','0','0','0','0','0','0',
        '0','0','0','0','0','0','0','0',
        '0','0','0','0','0','0','0','0',
        '0','0','0','0','0','0','0','0',
        -- *
        '0','0','0','0','0','0','0','0',
        '0','0','0','0','0','0','0','0',
        '0','0','0','0','0','0','0','0',
        '0','0','0','1','0','0','0','0',
        '0','1','0','1','0','1','0','0',
        '0','0','1','1','1','0','0','0',
        '0','0','1','0','1','0','0','0',
        '0','1','1','0','1','1','0','0',
        '0','0','1','0','1','0','0','0',
        '0','0','0','0','0','0','0','0',
        '0','0','0','0','0','0','0','0',
        '0','0','0','0','0','0','0','0',
        '0','0','0','0','0','0','0','0',
        '0','0','0','0','0','0','0','0',
        '0','0','0','0','0','0','0','0',
        '0','0','0','0','0','0','0','0',
        -- /
        '0','0','0','0','0','0','0','0',
        '0','0','0','0','0','0','0','0',
        '0','0','0','0','0','0','0','1',
        '0','0','0','0','0','0','1','0',
        '0','0','0','0','0','0','1','0',
        '0','0','0','0','0','0','1','0',
        '0','0','0','0','0','1','0','0',
        '0','0','0','0','0','1','0','0',
        '0','0','0','0','0','1','0','0',
        '0','0','0','0','1','0','0','0',
        '0','0','0','0','1','0','0','0',
        '0','0','0','0','1','0','0','0',
        '0','0','0','1','0','0','0','0',
        '0','0','0','1','0','0','0','0',
        '0','0','0','1','0','0','0','0',
        '0','0','1','0','0','0','0','0',
        --
        '0','0','0','0','0','0','0','0',
        '0','0','0','0','0','0','0','0',
        '0','0','0','0','0','0','0','0',
        '0','0','0','0','0','0','0','0',
        '0','0','0','0','0','0','0','0',
        '0','0','0','0','0','0','0','0',
        '0','0','0','0','0','0','0','0',
        '0','0','0','0','0','0','0','0',
        '0','0','0','0','0','0','0','0',
        '0','0','0','0','0','0','0','0',
        '0','0','0','0','0','0','0','0',
        '0','0','0','0','0','0','0','0',
        '0','0','0','0','0','0','0','0',
        '0','0','0','0','0','0','0','0',
        '0','0','0','0','0','0','0','0',
        '0','0','0','0','0','0','0','0'
        );
begin

    -- Clock divisor
    -- Divide system clock (100 MHz) by 4
    process(clk)
    begin
        if rising_edge(clk) then
            if rst='1' then
                ClkDiv <= (others => '0');
            else
                ClkDiv <= ClkDiv + 1;
            end if;
        end if;
    end process;

    -- 25 MHz clock (one system clock pulse width)
    Clk25 <= '1' when (ClkDiv = 3) else '0';


    -- Horizontal pixel counter

    process(clk)
    begin
        if rising_edge(clk) then
            if rst = '1' then
                Xpixel <= "0000000000";
            elsif Clk25='1' then
                if Xpixel = 799 then
                    Xpixel <= "0000000000";
                else
                    Xpixel <= Xpixel + 1;
                end if;
            end if;
        end if;
    end process;


    -- Horizontal sync

    -- ***********************************
    -- *                                 *
    -- *  VHDL for :                     *
    -- *  Hsync                          *
    -- *                                 *
    -- ***********************************

    process(Xpixel)
    begin
        if Xpixel>656 and Xpixel <=752 then
            Hsync<='0';
        else
            Hsync<='1';
        end if;
    end process;





    -- Vertical pixel counter

    -- ***********************************
    -- *                                 *
    -- *  VHDL for :                     *
    -- *  Ypixel                         *
    -- *                                 *
    -- ***********************************
    process(clk)
    begin
        if rising_edge(clk) then
            if rst='1' then
                Ypixel <= "0000000000";
            elsif Xpixel = 0 then
                if Ypixel = 520 then
                    Ypixel <= "0000000000";
                elsif Clk25='1' then
                    Ypixel <= Ypixel + 1;
                end if;
            end if;
        end if;
    end process;


    -- Vertical sync

    -- ***********************************
    -- *                                 *
    -- *  VHDL for :                     *
    -- *  Vsync                          *
    -- *                                 *
    -- ***********************************

    process(Ypixel)
    begin
        if Ypixel>490 and Ypixel <=492 then
            Vsync<='0';
        else
            Vsync<='1';
        end if;
    end process;

    -- Video blanking signal

    -- ***********************************
    -- *                                 *
    -- *  VHDL for :                     *
    -- *  Blank                          *
    -- *                                 *
    -- ***********************************
    process(Xpixel, Ypixel)
    begin
        if Ypixel >= 480 or Xpixel >= 640 then
            blank<='1';
        else
            blank<='0';
        end if;
    end process;
    --blank <= '1' when Ypixel > 480 and Xpixel > 640 else '0';




    -- Tile memory
    process(clk)
    begin
        if rising_edge(clk) then
            if (blank = '0') then
        		if tileRow = '1' and Xpixel>320 then
        		   tilepixel <= x"00";
                elsif Xpixel>320 then
        			tilepixel <= x"ff";
                elsif bitmem_in='1' then
                    tilepixel<=x"ff";
                else
                    tilepixel <= x"00";
        		end if;

                tileRow <= tileMem(to_integer(tileAddr));
            else
       		    tilePixel <= (others => '0');
                tileRow <= '0';
            end if;
        end if;
    end process;


    --with tileRow select tilePixel <=
      --  x"00" when '1',
      --  x"ff" when others;
   --tilepixel <= x"00";
    -- Tile memory address composite
    --tilecontent <= ;
    tileAddr <= unsigned(picmem_in(7 downto 0)) & Ypixel(3 downto 0) & Xpixel(2 downto 0);


    -- Picture memory address composite
    addr <= to_unsigned(80, 8) * Ypixel(8 downto 4) + Xpixel(9 downto 3);


    -- VGA generation
    vgaRed(2)   <= tilePixel(7);
    vgaRed(1)   <= tilePixel(6);
    vgaRed(0)   <= tilePixel(5);
    vgaGreen(2) <= tilePixel(4);
    vgaGreen(1) <= tilePixel(3);
    vgaGreen(0) <= tilePixel(2);
    vgaBlue(2)  <= tilePixel(1);
    vgaBlue(1)  <= tilePixel(0);


end Behavioral;

