--------------------------------------------------------------------------------
-- VGA MOTOR
-- Anders Nilsson
-- 16-feb-2016
-- Version 1.1


-- library declaration
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;            -- basic IEEE library
use IEEE.NUMERIC_STD.ALL;               -- IEEE library for the unsigned type


-- entity
entity VGA_MOTOR is
    port ( clk	  : in std_logic;
    	 data     : in std_logic_vector(7 downto 0);
    	 addr     : out unsigned(12 downto 0);
    	 rst      : in std_logic;
    	 vgaRed   : out std_logic_vector(2 downto 0);
    	 vgaGreen : out std_logic_vector(2 downto 0);
    	 vgaBlue  : out std_logic_vector(2 downto 1);
    	 Hsync    : out std_logic;
    	 Vsync    : out std_logic);
end VGA_MOTOR;


-- architecture
architecture Behavioral of VGA_MOTOR is

    signal Xpixel : unsigned(9 downto 0);         -- Horizontal pixel counter
    signal Ypixel : unsigned(9 downto 0);		-- Vertical pixel counter
    signal ClkDiv : unsigned(1 downto 0);		-- Clock divisor, to generate 25 MHz signal
    signal Clk25  : std_logic;			-- One pulse width 25 MHz signal

    signal tilePixel : std_logic_vector(7 downto 0);	-- Tile pixel data
    signal tileAddr  : unsigned(14 downto 0);	-- Tile address

    signal blank : std_logic;                    -- blanking signal
    signal tilerow : std_logic_vector(7 downto 0);

    -- Tile memory type
    type ram_t is array (0 to 767) of std_logic_vector(7 downto 0);

    -- Tile memory
    signal tileMem : ram_t :=(
    --
			"00000000",
			"00000000",
			"00000000",
			"00000000",
			"00000000",
			"00000000",
			"00000000",
			"00000000",
			"00000000",
			"00000000",
			"00000000",
			"00000000",
			"00000000",
			"00000000",
			"00000000",
			"00000000",
			-- A
			"00000000",
			"00000000",
			"00000000",
			"00010000",
			"00101000",
			"00101000",
			"00101000",
			"01000100",
			"01000100",
			"01111100",
			"01000100",
			"10000010",
			"10000010",
			"00000000",
			"00000000",
			"00000000",
			-- B
			"00000000",
			"00000000",
			"00000000",
			"01111100",
			"01000010",
			"01000010",
			"01000010",
			"01111100",
			"01000010",
			"01000010",
			"01000010",
			"01000010",
			"01111100",
			"00000000",
			"00000000",
			"00000000",
			-- C
			"00000000",
			"00000000",
			"00000000",
			"00011100",
			"00100010",
			"01000000",
			"01000000",
			"01000000",
			"01000000",
			"01000000",
			"01000000",
			"00100010",
			"00011100",
			"00000000",
			"00000000",
			"00000000",
			-- D
			"00000000",
			"00000000",
			"00000000",
			"01111000",
			"01000100",
			"01000010",
			"01000010",
			"01000010",
			"01000010",
			"01000010",
			"01000010",
			"01000100",
			"01111000",
			"00000000",
			"00000000",
			"00000000",
			-- E
			"00000000",
			"00000000",
			"00000000",
			"00111111",
			"00100000",
			"00100000",
			"00100000",
			"00111110",
			"00100000",
			"00100000",
			"00100000",
			"00100000",
			"00111111",
			"00000000",
			"00000000",
			"00000000",
			-- F
			"00000000",
			"00000000",
			"00000000",
			"00111111",
			"00100000",
			"00100000",
			"00100000",
			"00111110",
			"00100000",
			"00100000",
			"00100000",
			"00100000",
			"00100000",
			"00000000",
			"00000000",
			"00000000",
			-- G
			"00000000",
			"00000000",
			"00000000",
			"00011100",
			"00100010",
			"01000000",
			"01000000",
			"01000000",
			"01000010",
			"01000010",
			"01000010",
			"00100010",
			"00011110",
			"00000000",
			"00000000",
			"00000000",
			-- H
			"00000000",
			"00000000",
			"00000000",
			"01000010",
			"01000010",
			"01000010",
			"01000010",
			"01111110",
			"01000010",
			"01000010",
			"01000010",
			"01000010",
			"01000010",
			"00000000",
			"00000000",
			"00000000",
			-- I
			"00000000",
			"00000000",
			"00000000",
			"00111110",
			"00001000",
			"00001000",
			"00001000",
			"00001000",
			"00001000",
			"00001000",
			"00001000",
			"00001000",
			"00111110",
			"00000000",
			"00000000",
			"00000000",
			-- J
			"00000000",
			"00000000",
			"00000000",
			"00111110",
			"00000010",
			"00000010",
			"00000010",
			"00000010",
			"00000010",
			"00000010",
			"00000010",
			"01000010",
			"00111100",
			"00000000",
			"00000000",
			"00000000",
			-- K
			"00000000",
			"00000000",
			"00000000",
			"00100001",
			"00100010",
			"00100100",
			"00101000",
			"00110000",
			"00101000",
			"00100100",
			"00100100",
			"00100010",
			"00100001",
			"00000000",
			"00000000",
			"00000000",
			-- L
			"00000000",
			"00000000",
			"00000000",
			"00100000",
			"00100000",
			"00100000",
			"00100000",
			"00100000",
			"00100000",
			"00100000",
			"00100000",
			"00100000",
			"00111111",
			"00000000",
			"00000000",
			"00000000",
			-- M
			"00000000",
			"00000000",
			"00000000",
			"00100100",
			"00100100",
			"00100100",
			"01011010",
			"01011010",
			"01011010",
			"01000010",
			"01000010",
			"01000010",
			"01000010",
			"00000000",
			"00000000",
			"00000000",
			-- N
			"00000000",
			"00000000",
			"00000000",
			"01000010",
			"01100010",
			"01100010",
			"01010010",
			"01011010",
			"01001010",
			"01001010",
			"01000110",
			"01000110",
			"01000010",
			"00000000",
			"00000000",
			"00000000",
			-- O
			"00000000",
			"00000000",
			"00000000",
			"00011000",
			"00100100",
			"01000010",
			"01000010",
			"01000010",
			"01000010",
			"01000010",
			"01000010",
			"00100100",
			"00011000",
			"00000000",
			"00000000",
			"00000000",
			-- P
			"00000000",
			"00000000",
			"00000000",
			"00111110",
			"00100001",
			"00100001",
			"00100001",
			"00100001",
			"00111110",
			"00100000",
			"00100000",
			"00100000",
			"00100000",
			"00000000",
			"00000000",
			"00000000",
			-- Q
			"00000000",
			"00000000",
			"00000000",
			"00011000",
			"00100100",
			"01000010",
			"01000010",
			"01000010",
			"01000010",
			"01000010",
			"01000010",
			"00100100",
			"00011000",
			"00011000",
			"00000110",
			"00000000",
			-- R
			"00000000",
			"00000000",
			"00000000",
			"01111100",
			"01000010",
			"01000010",
			"01000010",
			"01000010",
			"01111100",
			"01001000",
			"01000100",
			"01000010",
			"01000001",
			"00000000",
			"00000000",
			"00000000",
			-- S
			"00000000",
			"00000000",
			"00000000",
			"00111100",
			"01000010",
			"01000000",
			"01000000",
			"00110000",
			"00001100",
			"00000010",
			"00000010",
			"01000010",
			"01111100",
			"00000000",
			"00000000",
			"00000000",
			-- T
			"00000000",
			"00000000",
			"00000000",
			"11111110",
			"00010000",
			"00010000",
			"00010000",
			"00010000",
			"00010000",
			"00010000",
			"00010000",
			"00010000",
			"00010000",
			"00000000",
			"00000000",
			"00000000",
			-- U
			"00000000",
			"00000000",
			"00000000",
			"01000010",
			"01000010",
			"01000010",
			"01000010",
			"01000010",
			"01000010",
			"01000010",
			"01000010",
			"01000010",
			"00111100",
			"00000000",
			"00000000",
			"00000000",
			-- V
			"00000000",
			"00000000",
			"00000000",
			"10000010",
			"10000010",
			"01000100",
			"01000100",
			"01000100",
			"01100100",
			"00101000",
			"00101000",
			"00111000",
			"00010000",
			"00000000",
			"00000000",
			"00000000",
			-- W
			"00000000",
			"00000000",
			"00000000",
			"01000010",
			"01000010",
			"01000010",
			"01000010",
			"01011010",
			"01011010",
			"01011010",
			"01100110",
			"01100110",
			"01000010",
			"00000000",
			"00000000",
			"00000000",
			-- X
			"00000000",
			"00000000",
			"00000000",
			"10000010",
			"01000100",
			"01000100",
			"00101000",
			"00010000",
			"00010000",
			"00101000",
			"01000100",
			"01000100",
			"10000010",
			"00000000",
			"00000000",
			"00000000",
			-- Y
			"00000000",
			"00000000",
			"00000000",
			"10000010",
			"01000100",
			"01000100",
			"00101000",
			"00101000",
			"00010000",
			"00010000",
			"00010000",
			"00010000",
			"00010000",
			"00000000",
			"00000000",
			"00000000",
			-- Z
			"00000000",
			"00000000",
			"00000000",
			"01111110",
			"00000010",
			"00000100",
			"00001000",
			"00001000",
			"00010000",
			"00110000",
			"00100000",
			"01000000",
			"01111110",
			"00000000",
			"00000000",
			"00000000",
			-- Å
			"00011000",
			"00100100",
			"00100100",
			"00011000",
			"00011000",
			"00100100",
			"00100100",
			"00100100",
			"01000010",
			"01111110",
			"01000010",
			"10000011",
			"10000001",
			"00000000",
			"00000000",
			"00000000",
			-- Ä
			"00101000",
			"00101000",
			"00000000",
			"00010000",
			"00101000",
			"00101000",
			"00101000",
			"01000100",
			"01000100",
			"01111100",
			"01000100",
			"10000010",
			"10000010",
			"00000000",
			"00000000",
			"00000000",
			-- Ö
			"00010100",
			"00010100",
			"00000000",
			"00011000",
			"00100100",
			"01000010",
			"01000010",
			"01000010",
			"01000010",
			"01000010",
			"01000010",
			"00100100",
			"00011000",
			"00000000",
			"00000000",
			"00000000",
			-- 1
			"00000000",
			"00000000",
			"00000000",
			"00000100",
			"00001100",
			"00010100",
			"00000100",
			"00000100",
			"00000100",
			"00000100",
			"00000100",
			"00000100",
			"00011111",
			"00000000",
			"00000000",
			"00000000",
			-- 2
			"00000000",
			"00000000",
			"00000000",
			"00111100",
			"01000010",
			"00000010",
			"00000010",
			"00000100",
			"00001000",
			"00010000",
			"00100000",
			"01000000",
			"01111110",
			"00000000",
			"00000000",
			"00000000",
			-- 3
			"00000000",
			"00000000",
			"00000000",
			"01111100",
			"00000010",
			"00000010",
			"00000010",
			"00011100",
			"00000010",
			"00000010",
			"00000010",
			"00000010",
			"01111100",
			"00000000",
			"00000000",
			"00000000",
			-- 4
			"00000000",
			"00000000",
			"00000000",
			"00000100",
			"00001100",
			"00010100",
			"00100100",
			"00100100",
			"01000100",
			"01111110",
			"00000100",
			"00000100",
			"00000100",
			"00000000",
			"00000000",
			"00000000",
			-- 5
			"00000000",
			"00000000",
			"00000000",
			"00011111",
			"00010000",
			"00010000",
			"00010000",
			"00011100",
			"00000010",
			"00000001",
			"00000001",
			"00000010",
			"00111100",
			"00000000",
			"00000000",
			"00000000",
			-- 6
			"00000000",
			"00000000",
			"00000000",
			"00001100",
			"00010000",
			"00100000",
			"01000000",
			"01111100",
			"01000010",
			"01000010",
			"01000010",
			"00100100",
			"00011000",
			"00000000",
			"00000000",
			"00000000",
			-- 7
			"00000000",
			"00000000",
			"00000000",
			"00111111",
			"00000001",
			"00000010",
			"00000100",
			"00000100",
			"00001000",
			"00001000",
			"00010000",
			"00010000",
			"00010000",
			"00000000",
			"00000000",
			"00000000",
			-- 8
			"00000000",
			"00000000",
			"00000000",
			"00111100",
			"01000010",
			"01000010",
			"01000010",
			"00111100",
			"00101100",
			"01000010",
			"01000010",
			"01000010",
			"00111100",
			"00000000",
			"00000000",
			"00000000",
			-- 9
			"00000000",
			"00000000",
			"00000000",
			"00111000",
			"01000100",
			"01000010",
			"01000010",
			"01000010",
			"00111110",
			"00000010",
			"00000100",
			"00001000",
			"00110000",
			"00000000",
			"00000000",
			"00000000",
			-- 0
			"00000000",
			"00000000",
			"00000000",
			"00011000",
			"00100100",
			"01000010",
			"01000010",
			"01011010",
			"01011010",
			"01000010",
			"01000010",
			"00100100",
			"00011000",
			"00000000",
			"00000000",
			"00000000",
			-- π
			"00000000",
			"00000000",
			"00000000",
			"00000000",
			"00000000",
			"00000000",
			"00111111",
			"00100001",
			"00100001",
			"00100001",
			"00100001",
			"00100001",
			"00100001",
			"00000000",
			"00000000",
			"00000000",
			-- Ω
			"00000000",
			"00000000",
			"00000000",
			"00011000",
			"00100100",
			"01000010",
			"01000010",
			"01000010",
			"01000010",
			"01000010",
			"01000010",
			"00100100",
			"01100110",
			"00000000",
			"00000000",
			"00000000",
			-- .
			"00000000",
			"00000000",
			"00000000",
			"00000000",
			"00000000",
			"00000000",
			"00000000",
			"00000000",
			"00000000",
			"00000000",
			"00000000",
			"00000000",
			"00001000",
			"00000000",
			"00000000",
			"00000000",
			-- =
			"00000000",
			"00000000",
			"00000000",
			"00000000",
			"00000000",
			"00000000",
			"00000000",
			"01111110",
			"00000000",
			"00000000",
			"01111110",
			"00000000",
			"00000000",
			"00000000",
			"00000000",
			"00000000",
			-- +
			"00000000",
			"00000000",
			"00000000",
			"00000000",
			"00000000",
			"00010000",
			"00010000",
			"00010000",
			"11111110",
			"00010000",
			"00010000",
			"00010000",
			"00000000",
			"00000000",
			"00000000",
			"00000000",
			-- -
			"00000000",
			"00000000",
			"00000000",
			"00000000",
			"00000000",
			"00000000",
			"00000000",
			"00000000",
			"00000000",
			"00011110",
			"00000000",
			"00000000",
			"00000000",
			"00000000",
			"00000000",
			"00000000",
			-- *
			"00000000",
			"00000000",
			"00000000",
			"00010000",
			"01010100",
			"00111000",
			"00101000",
			"01101100",
			"00101000",
			"00000000",
			"00000000",
			"00000000",
			"00000000",
			"00000000",
			"00000000",
			"00000000",
			-- /
			"00000000",
			"00000000",
			"00000001",
			"00000010",
			"00000010",
			"00000010",
			"00000100",
			"00000100",
			"00000100",
			"00001000",
			"00001000",
			"00001000",
			"00010000",
			"00010000",
			"00010000",
			"00100000"
                );

begin

    -- Clock divisor
    -- Divide system clock (100 MHz) by 4
    process(clk)
    begin
        if rising_edge(clk) then
            if rst='1' then
                ClkDiv <= (others => '0');
            else
                ClkDiv <= ClkDiv + 1;
            end if;
        end if;
    end process;

    -- 25 MHz clock (one system clock pulse width)
    Clk25 <= '1' when (ClkDiv = 3) else '0';


    -- Horizontal pixel counter

    process(clk)
    begin
        if rising_edge(clk) then
            if rst = '1' then
                Xpixel <= "0000000000";
            elsif Clk25='1' then
                if Xpixel = 799 then
                    Xpixel <= "0000000000";
                else
                    Xpixel <= Xpixel + 1;
                end if;
            end if;
        end if;
    end process;


    -- Horizontal sync

    -- ***********************************
    -- *                                 *
    -- *  VHDL for :                     *
    -- *  Hsync                          *
    -- *                                 *
    -- ***********************************

    process(Xpixel)
    begin
        if Xpixel>656 and Xpixel <=752 then
            Hsync<='0';
        else
            Hsync<='1';
        end if;
    end process;





    -- Vertical pixel counter

    -- ***********************************
    -- *                                 *
    -- *  VHDL for :                     *
    -- *  Ypixel                         *
    -- *                                 *
    -- ***********************************
    process(clk)
    begin
        if rising_edge(clk) then
            if rst='1' then
                Ypixel <= "0000000000";
            elsif Xpixel = 0 then
                if Ypixel = 520 then
                    Ypixel <= "0000000000";
                elsif Clk25='1' then
                    Ypixel <= Ypixel + 1;
                end if;
            end if;
        end if;
    end process;


    -- Vertical sync

    -- ***********************************
    -- *                                 *
    -- *  VHDL for :                     *
    -- *  Vsync                          *
    -- *                                 *
    -- ***********************************

    process(Ypixel)
    begin
        if Ypixel>490 and Ypixel <=492 then
            Vsync<='0';
        else
            Vsync<='1';
        end if;
    end process;

    -- Video blanking signal

    -- ***********************************
    -- *                                 *
    -- *  VHDL for :                     *
    -- *  Blank                          *
    -- *                                 *
    -- ***********************************
    process(Xpixel, Ypixel)
    begin
        if Ypixel >= 480 or Xpixel >= 640 then
            blank<='1';
        else
            blank<='0';
        end if;
    end process;
    --blank <= '1' when Ypixel > 480 and Xpixel > 640 else '0';




    -- Tile memory
    process(clk)
    begin
        if rising_edge(clk) then
            if (blank = '0') then
                tileRow <= tilemem(to_integer(unsigned(data)*16+unsigned(Ypixel(3 downto 0))));
            else
                tileRow <= (others => '0');
            end if;
        end if;
    end process;


    -- TODO: Probaly off by one char
    process(clk)
    begin
        if rising_edge(clk) then
            if tileRow(to_integer(Xpixel(2 downto 0)))='1' then
                tilePixel <= x"00";
            else
                tilePixel <= x"ff";
            end if;
        end if;
    end process;
    -- Tile memory address composite
    --tilecontent <= ;
    tileAddr <= unsigned(data(7 downto 0)) & Ypixel(3 downto 0) & Xpixel(2 downto 0);


    -- Picture memory address composite
    addr <= to_unsigned(40, 8) * Ypixel(8 downto 4) + Xpixel(9 downto 3);


    -- VGA generation
    vgaRed(2)   <= tilePixel(7);
    vgaRed(1)   <= tilePixel(6);
    vgaRed(0)   <= tilePixel(5);
    vgaGreen(2) <= tilePixel(4);
    vgaGreen(1) <= tilePixel(3);
    vgaGreen(0) <= tilePixel(2);
    vgaBlue(2)  <= tilePixel(1);
    vgaBlue(1)  <= tilePixel(0);


end Behavioral;
